----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    02:40:04 07/01/2022 
-- Design Name: 
-- Module Name:    DFF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lsfit2_model is

Port ( clk,nrst,enb,D : in  STD_LOGIC;
             Q,nQ: out std_logic);

end lsfit2_model;

architecture Behavioral of lsfit2_model is

begin
process(clk,enb,D,nrst)
begin
	if(enb ='0')then
		Q <= 'Z';
		nQ <= 'Z';
		elsif (nrst = '1') then
			Q <= '0';
			nQ <= '1';
			elsif(clk'event and clk ='1') then
			Q <= D;
			nQ <= not D;
			end if;
end process;

end Behavioral;

